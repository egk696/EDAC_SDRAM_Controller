OBUF_inst : OBUF PORT MAP (
		datain	 => datain_sig,
		dataout	 => dataout_sig
	);
