-- EDAC_SDRAM_Controller_Demo.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity EDAC_SDRAM_Controller_Demo is
	port (
		debug_err_counter_o        : out   std_logic_vector(31 downto 0);                    --        debug.err_counter_o
		debug_err_detect_o         : out   std_logic;                                        --             .err_detect_o
		debug_healing_proc_run_o   : out   std_logic;                                        --             .healing_proc_run_o
		debug_mem_ready_o          : out   std_logic;                                        --             .mem_ready_o
		debug_scrubbing_proc_run_o : out   std_logic;                                        --             .scrubbing_proc_run_o
		debug_voted_data_o         : out   std_logic_vector(31 downto 0);                    --             .voted_data_o
		sdram_cke_o                : out   std_logic;                                        --        sdram.cke_o
		sdram_bank_o               : out   std_logic_vector(1 downto 0);                     --             .bank_o
		sdram_addr_o               : out   std_logic_vector(12 downto 0);                    --             .addr_o
		sdram_cs_o                 : out   std_logic;                                        --             .cs_o
		sdram_ras_o                : out   std_logic;                                        --             .ras_o
		sdram_cas_o                : out   std_logic;                                        --             .cas_o
		sdram_we_o                 : out   std_logic;                                        --             .we_o
		sdram_dqm_o                : out   std_logic_vector(3 downto 0);                     --             .dqm_o
		sdram_dataQ_io             : inout std_logic_vector(31 downto 0) := (others => '0'); --             .dataQ_io
		sevensegment_hex7          : out   std_logic_vector(6 downto 0);                     -- sevensegment.hex7
		sevensegment_hex6          : out   std_logic_vector(6 downto 0);                     --             .hex6
		sevensegment_hex5          : out   std_logic_vector(6 downto 0);                     --             .hex5
		sevensegment_hex4          : out   std_logic_vector(6 downto 0);                     --             .hex4
		sevensegment_hex3          : out   std_logic_vector(6 downto 0);                     --             .hex3
		sevensegment_hex2          : out   std_logic_vector(6 downto 0);                     --             .hex2
		sevensegment_hex1          : out   std_logic_vector(6 downto 0);                     --             .hex1
		sevensegment_hex0          : out   std_logic_vector(6 downto 0);                     --             .hex0
		sys_clk_clk                : in    std_logic                     := '0';             --      sys_clk.clk
		sys_rst_reset_n            : in    std_logic                     := '0'              --      sys_rst.reset_n
	);
end entity EDAC_SDRAM_Controller_Demo;

architecture rtl of EDAC_SDRAM_Controller_Demo is
	component sdram_ctrl_tmr_avs_multiport_interface is
		generic (
			DATA_WIDTH           : integer := 32;
			DQM_WIDTH            : integer := 2;
			ROW_WIDTH            : integer := 13;
			COLS_WIDTH           : integer := 10;
			BANK_WIDTH           : integer := 2;
			NOP_BOOT_CYCLES      : integer := 10000;
			REF_PERIOD           : integer := 92;
			REF_COMMAND_COUNT    : integer := 8;
			REF_COMMAND_PERIOD   : integer := 8;
			PRECH_COMMAND_PERIOD : integer := 2;
			ACT_TO_RW_CYCLES     : integer := 2;
			IN_DATA_TO_PRE       : integer := 2;
			CAS_LAT_CYCLES       : integer := 2;
			MODE_REG_CYCLES      : integer := 2;
			BURST_LENGTH         : integer := 0;
			DRIVE_STRENGTH       : integer := 0;
			RAM_COLS             : integer := 1024;
			RAM_ROWS             : integer := 8192;
			RAM_BANKS            : integer := 4;
			TMR_COLS             : integer := 768;
			SCRUBBER_WAIT_CYCLES : integer := 64;
			EXT_MODE_REG_EN      : boolean := true;
			GEN_ERR_INJ          : boolean := false
		);
		port (
			rsi_reset_n          : in    std_logic                     := 'X';             -- reset_n
			portA_address        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			portA_read           : in    std_logic                     := 'X';             -- read
			portA_readdata       : out   std_logic_vector(31 downto 0);                    -- readdata
			portA_write          : in    std_logic                     := 'X';             -- write
			portA_writedata      : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			portA_waitrequest    : out   std_logic;                                        -- waitrequest
			portA_readdatavalid  : out   std_logic;                                        -- readdatavalid
			portB_address        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			portB_read           : in    std_logic                     := 'X';             -- read
			portB_readdata       : out   std_logic_vector(31 downto 0);                    -- readdata
			portB_write          : in    std_logic                     := 'X';             -- write
			portB_writedata      : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			portB_waitrequest    : out   std_logic;                                        -- waitrequest
			portB_readdatavalid  : out   std_logic;                                        -- readdatavalid
			csi_clock            : in    std_logic                     := 'X';             -- clk
			err_counter_o        : out   std_logic_vector(31 downto 0);                    -- err_counter_o
			err_detect_o         : out   std_logic;                                        -- err_detect_o
			healing_proc_run_o   : out   std_logic;                                        -- healing_proc_run_o
			mem_ready_o          : out   std_logic;                                        -- mem_ready_o
			scrubbing_proc_run_o : out   std_logic;                                        -- scrubbing_proc_run_o
			voted_data_o         : out   std_logic_vector(31 downto 0);                    -- voted_data_o
			cke_o                : out   std_logic;                                        -- cke_o
			bank_o               : out   std_logic_vector(1 downto 0);                     -- bank_o
			addr_o               : out   std_logic_vector(12 downto 0);                    -- addr_o
			cs_o                 : out   std_logic;                                        -- cs_o
			ras_o                : out   std_logic;                                        -- ras_o
			cas_o                : out   std_logic;                                        -- cas_o
			we_o                 : out   std_logic;                                        -- we_o
			dqm_o                : out   std_logic_vector(3 downto 0);                     -- dqm_o
			dataQ_io             : inout std_logic_vector(31 downto 0) := (others => 'X')  -- dataQ_io
		);
	end component sdram_ctrl_tmr_avs_multiport_interface;

	component EDAC_SDRAM_Controller_Demo_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(27 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(27 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component EDAC_SDRAM_Controller_Demo_nios2_gen2_0;

	component EDAC_SDRAM_Controller_Demo_onchip_memory2_0 is
		port (
			address     : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			address2    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk         : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			freeze      : in  std_logic                     := 'X'              -- freeze
		);
	end component EDAC_SDRAM_Controller_Demo_onchip_memory2_0;

	component sevensegment_avalon_master_interface is
		generic (
			DATA_WIDTH    : integer := 32;
			ADDRESS_WIDTH : integer := 25;
			UPDATE_RATE   : integer := 128
		);
		port (
			avm_address       : out std_logic_vector(24 downto 0);                    -- address
			avm_read          : out std_logic;                                        -- read
			avm_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avm_write         : out std_logic;                                        -- write
			avm_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			avm_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			avm_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			rsi_reset_n       : in  std_logic                     := 'X';             -- reset_n
			HEX7              : out std_logic_vector(6 downto 0);                     -- hex7
			HEX6              : out std_logic_vector(6 downto 0);                     -- hex6
			HEX5              : out std_logic_vector(6 downto 0);                     -- hex5
			HEX4              : out std_logic_vector(6 downto 0);                     -- hex4
			HEX3              : out std_logic_vector(6 downto 0);                     -- hex3
			HEX2              : out std_logic_vector(6 downto 0);                     -- hex2
			HEX1              : out std_logic_vector(6 downto 0);                     -- hex1
			HEX0              : out std_logic_vector(6 downto 0);                     -- hex0
			csi_clock         : in  std_logic                     := 'X'              -- clk
		);
	end component sevensegment_avalon_master_interface;

	component EDAC_SDRAM_Controller_Demo_mm_interconnect_1 is
		port (
			clk_0_clk_clk                                  : in  std_logic                     := 'X';             -- clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_data_master_address               : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest           : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                  : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_write                 : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address        : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read           : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			edac_sdram_controller_0_porta_address          : out std_logic_vector(24 downto 0);                    -- address
			edac_sdram_controller_0_porta_write            : out std_logic;                                        -- write
			edac_sdram_controller_0_porta_read             : out std_logic;                                        -- read
			edac_sdram_controller_0_porta_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			edac_sdram_controller_0_porta_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			edac_sdram_controller_0_porta_readdatavalid    : in  std_logic                     := 'X';             -- readdatavalid
			edac_sdram_controller_0_porta_waitrequest      : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write             : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read              : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
			onchip_memory2_0_s1_address                    : out std_logic_vector(12 downto 0);                    -- address
			onchip_memory2_0_s1_write                      : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                 : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                 : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                      : out std_logic;                                        -- clken
			onchip_memory2_0_s2_address                    : out std_logic_vector(12 downto 0);                    -- address
			onchip_memory2_0_s2_write                      : out std_logic;                                        -- write
			onchip_memory2_0_s2_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s2_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s2_byteenable                 : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s2_chipselect                 : out std_logic;                                        -- chipselect
			onchip_memory2_0_s2_clken                      : out std_logic                                         -- clken
		);
	end component EDAC_SDRAM_Controller_Demo_mm_interconnect_1;

	component EDAC_SDRAM_Controller_Demo_irq_mapper is
		port (
			clk        : in  std_logic                     := 'X'; -- clk
			reset      : in  std_logic                     := 'X'; -- reset
			sender_irq : out std_logic_vector(31 downto 0)         -- irq
		);
	end component EDAC_SDRAM_Controller_Demo_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal sevensegment_avalon_master_interface_0_avalon_master_0_readdata      : std_logic_vector(31 downto 0); -- edac_sdram_controller_0:portB_readdata -> sevensegment_avalon_master_interface_0:avm_readdata
	signal sevensegment_avalon_master_interface_0_avalon_master_0_waitrequest   : std_logic;                     -- edac_sdram_controller_0:portB_waitrequest -> sevensegment_avalon_master_interface_0:avm_waitrequest
	signal sevensegment_avalon_master_interface_0_avalon_master_0_address       : std_logic_vector(24 downto 0); -- sevensegment_avalon_master_interface_0:avm_address -> edac_sdram_controller_0:portB_address
	signal sevensegment_avalon_master_interface_0_avalon_master_0_read          : std_logic;                     -- sevensegment_avalon_master_interface_0:avm_read -> edac_sdram_controller_0:portB_read
	signal sevensegment_avalon_master_interface_0_avalon_master_0_readdatavalid : std_logic;                     -- edac_sdram_controller_0:portB_readdatavalid -> sevensegment_avalon_master_interface_0:avm_readdatavalid
	signal sevensegment_avalon_master_interface_0_avalon_master_0_write         : std_logic;                     -- sevensegment_avalon_master_interface_0:avm_write -> edac_sdram_controller_0:portB_write
	signal sevensegment_avalon_master_interface_0_avalon_master_0_writedata     : std_logic_vector(31 downto 0); -- sevensegment_avalon_master_interface_0:avm_writedata -> edac_sdram_controller_0:portB_writedata
	signal nios2_gen2_0_data_master_readdata                                    : std_logic_vector(31 downto 0); -- mm_interconnect_1:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                                 : std_logic;                     -- mm_interconnect_1:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                                 : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_1:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                     : std_logic_vector(27 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_1:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                                  : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_1:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                        : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_1:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_write                                       : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_1:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                                   : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_1:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                             : std_logic_vector(31 downto 0); -- mm_interconnect_1:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                          : std_logic;                     -- mm_interconnect_1:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                              : std_logic_vector(27 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_1:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                                 : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_1:nios2_gen2_0_instruction_master_read
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata              : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_1:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest           : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_1:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess           : std_logic;                     -- mm_interconnect_1:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address               : std_logic_vector(8 downto 0);  -- mm_interconnect_1:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read                  : std_logic;                     -- mm_interconnect_1:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable            : std_logic_vector(3 downto 0);  -- mm_interconnect_1:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write                 : std_logic;                     -- mm_interconnect_1:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_1:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_1_edac_sdram_controller_0_porta_readdata             : std_logic_vector(31 downto 0); -- edac_sdram_controller_0:portA_readdata -> mm_interconnect_1:edac_sdram_controller_0_porta_readdata
	signal mm_interconnect_1_edac_sdram_controller_0_porta_waitrequest          : std_logic;                     -- edac_sdram_controller_0:portA_waitrequest -> mm_interconnect_1:edac_sdram_controller_0_porta_waitrequest
	signal mm_interconnect_1_edac_sdram_controller_0_porta_address              : std_logic_vector(24 downto 0); -- mm_interconnect_1:edac_sdram_controller_0_porta_address -> edac_sdram_controller_0:portA_address
	signal mm_interconnect_1_edac_sdram_controller_0_porta_read                 : std_logic;                     -- mm_interconnect_1:edac_sdram_controller_0_porta_read -> edac_sdram_controller_0:portA_read
	signal mm_interconnect_1_edac_sdram_controller_0_porta_readdatavalid        : std_logic;                     -- edac_sdram_controller_0:portA_readdatavalid -> mm_interconnect_1:edac_sdram_controller_0_porta_readdatavalid
	signal mm_interconnect_1_edac_sdram_controller_0_porta_write                : std_logic;                     -- mm_interconnect_1:edac_sdram_controller_0_porta_write -> edac_sdram_controller_0:portA_write
	signal mm_interconnect_1_edac_sdram_controller_0_porta_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_1:edac_sdram_controller_0_porta_writedata -> edac_sdram_controller_0:portA_writedata
	signal mm_interconnect_1_onchip_memory2_0_s1_chipselect                     : std_logic;                     -- mm_interconnect_1:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_1_onchip_memory2_0_s1_readdata                       : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_1:onchip_memory2_0_s1_readdata
	signal mm_interconnect_1_onchip_memory2_0_s1_address                        : std_logic_vector(12 downto 0); -- mm_interconnect_1:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_1_onchip_memory2_0_s1_byteenable                     : std_logic_vector(3 downto 0);  -- mm_interconnect_1:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_1_onchip_memory2_0_s1_write                          : std_logic;                     -- mm_interconnect_1:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_1_onchip_memory2_0_s1_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_1:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_1_onchip_memory2_0_s1_clken                          : std_logic;                     -- mm_interconnect_1:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal mm_interconnect_1_onchip_memory2_0_s2_chipselect                     : std_logic;                     -- mm_interconnect_1:onchip_memory2_0_s2_chipselect -> onchip_memory2_0:chipselect2
	signal mm_interconnect_1_onchip_memory2_0_s2_readdata                       : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata2 -> mm_interconnect_1:onchip_memory2_0_s2_readdata
	signal mm_interconnect_1_onchip_memory2_0_s2_address                        : std_logic_vector(12 downto 0); -- mm_interconnect_1:onchip_memory2_0_s2_address -> onchip_memory2_0:address2
	signal mm_interconnect_1_onchip_memory2_0_s2_byteenable                     : std_logic_vector(3 downto 0);  -- mm_interconnect_1:onchip_memory2_0_s2_byteenable -> onchip_memory2_0:byteenable2
	signal mm_interconnect_1_onchip_memory2_0_s2_write                          : std_logic;                     -- mm_interconnect_1:onchip_memory2_0_s2_write -> onchip_memory2_0:write2
	signal mm_interconnect_1_onchip_memory2_0_s2_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_1:onchip_memory2_0_s2_writedata -> onchip_memory2_0:writedata2
	signal mm_interconnect_1_onchip_memory2_0_s2_clken                          : std_logic;                     -- mm_interconnect_1:onchip_memory2_0_s2_clken -> onchip_memory2_0:clken2
	signal nios2_gen2_0_irq_irq                                                 : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal rst_controller_reset_out_reset                                       : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_1:nios2_gen2_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                   : std_logic;                     -- rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	signal sys_rst_reset_n_ports_inv                                            : std_logic;                     -- sys_rst_reset_n:inv -> rst_controller:reset_in0
	signal rst_controller_reset_out_reset_ports_inv                             : std_logic;                     -- rst_controller_reset_out_reset:inv -> [edac_sdram_controller_0:rsi_reset_n, nios2_gen2_0:reset_n, sevensegment_avalon_master_interface_0:rsi_reset_n]

begin

	edac_sdram_controller_0 : component sdram_ctrl_tmr_avs_multiport_interface
		generic map (
			DATA_WIDTH           => 32,
			DQM_WIDTH            => 4,
			ROW_WIDTH            => 13,
			COLS_WIDTH           => 10,
			BANK_WIDTH           => 2,
			NOP_BOOT_CYCLES      => 20000,
			REF_PERIOD           => 350,
			REF_COMMAND_COUNT    => 8,
			REF_COMMAND_PERIOD   => 8,
			PRECH_COMMAND_PERIOD => 2,
			ACT_TO_RW_CYCLES     => 2,
			IN_DATA_TO_PRE       => 2,
			CAS_LAT_CYCLES       => 2,
			MODE_REG_CYCLES      => 2,
			BURST_LENGTH         => 0,
			DRIVE_STRENGTH       => 0,
			RAM_COLS             => 1024,
			RAM_ROWS             => 8192,
			RAM_BANKS            => 4,
			TMR_COLS             => 768,
			SCRUBBER_WAIT_CYCLES => 64,
			EXT_MODE_REG_EN      => false,
			GEN_ERR_INJ          => false
		)
		port map (
			rsi_reset_n          => rst_controller_reset_out_reset_ports_inv,                             -- reset.reset_n
			portA_address        => mm_interconnect_1_edac_sdram_controller_0_porta_address,              -- porta.address
			portA_read           => mm_interconnect_1_edac_sdram_controller_0_porta_read,                 --      .read
			portA_readdata       => mm_interconnect_1_edac_sdram_controller_0_porta_readdata,             --      .readdata
			portA_write          => mm_interconnect_1_edac_sdram_controller_0_porta_write,                --      .write
			portA_writedata      => mm_interconnect_1_edac_sdram_controller_0_porta_writedata,            --      .writedata
			portA_waitrequest    => mm_interconnect_1_edac_sdram_controller_0_porta_waitrequest,          --      .waitrequest
			portA_readdatavalid  => mm_interconnect_1_edac_sdram_controller_0_porta_readdatavalid,        --      .readdatavalid
			portB_address        => sevensegment_avalon_master_interface_0_avalon_master_0_address,       -- portb.address
			portB_read           => sevensegment_avalon_master_interface_0_avalon_master_0_read,          --      .read
			portB_readdata       => sevensegment_avalon_master_interface_0_avalon_master_0_readdata,      --      .readdata
			portB_write          => sevensegment_avalon_master_interface_0_avalon_master_0_write,         --      .write
			portB_writedata      => sevensegment_avalon_master_interface_0_avalon_master_0_writedata,     --      .writedata
			portB_waitrequest    => sevensegment_avalon_master_interface_0_avalon_master_0_waitrequest,   --      .waitrequest
			portB_readdatavalid  => sevensegment_avalon_master_interface_0_avalon_master_0_readdatavalid, --      .readdatavalid
			csi_clock            => sys_clk_clk,                                                          -- clock.clk
			err_counter_o        => debug_err_counter_o,                                                  -- debug.err_counter_o
			err_detect_o         => debug_err_detect_o,                                                   --      .err_detect_o
			healing_proc_run_o   => debug_healing_proc_run_o,                                             --      .healing_proc_run_o
			mem_ready_o          => debug_mem_ready_o,                                                    --      .mem_ready_o
			scrubbing_proc_run_o => debug_scrubbing_proc_run_o,                                           --      .scrubbing_proc_run_o
			voted_data_o         => debug_voted_data_o,                                                   --      .voted_data_o
			cke_o                => sdram_cke_o,                                                          -- sdram.cke_o
			bank_o               => sdram_bank_o,                                                         --      .bank_o
			addr_o               => sdram_addr_o,                                                         --      .addr_o
			cs_o                 => sdram_cs_o,                                                           --      .cs_o
			ras_o                => sdram_ras_o,                                                          --      .ras_o
			cas_o                => sdram_cas_o,                                                          --      .cas_o
			we_o                 => sdram_we_o,                                                           --      .we_o
			dqm_o                => sdram_dqm_o,                                                          --      .dqm_o
			dataQ_io             => sdram_dataQ_io                                                        --      .dataQ_io
		);

	nios2_gen2_0 : component EDAC_SDRAM_Controller_Demo_nios2_gen2_0
		port map (
			clk                                 => sys_clk_clk,                                                --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                   --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                         --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                                       --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	onchip_memory2_0 : component EDAC_SDRAM_Controller_Demo_onchip_memory2_0
		port map (
			address     => mm_interconnect_1_onchip_memory2_0_s1_address,    --     s1.address
			clken       => mm_interconnect_1_onchip_memory2_0_s1_clken,      --       .clken
			chipselect  => mm_interconnect_1_onchip_memory2_0_s1_chipselect, --       .chipselect
			write       => mm_interconnect_1_onchip_memory2_0_s1_write,      --       .write
			readdata    => mm_interconnect_1_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_1_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_1_onchip_memory2_0_s1_byteenable, --       .byteenable
			address2    => mm_interconnect_1_onchip_memory2_0_s2_address,    --     s2.address
			chipselect2 => mm_interconnect_1_onchip_memory2_0_s2_chipselect, --       .chipselect
			clken2      => mm_interconnect_1_onchip_memory2_0_s2_clken,      --       .clken
			write2      => mm_interconnect_1_onchip_memory2_0_s2_write,      --       .write
			readdata2   => mm_interconnect_1_onchip_memory2_0_s2_readdata,   --       .readdata
			writedata2  => mm_interconnect_1_onchip_memory2_0_s2_writedata,  --       .writedata
			byteenable2 => mm_interconnect_1_onchip_memory2_0_s2_byteenable, --       .byteenable
			clk         => sys_clk_clk,                                      --   clk1.clk
			reset       => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,               --       .reset_req
			freeze      => '0'                                               -- (terminated)
		);

	sevensegment_avalon_master_interface_0 : component sevensegment_avalon_master_interface
		generic map (
			DATA_WIDTH    => 32,
			ADDRESS_WIDTH => 25,
			UPDATE_RATE   => 128
		)
		port map (
			avm_address       => sevensegment_avalon_master_interface_0_avalon_master_0_address,       --  avalon_master_0.address
			avm_read          => sevensegment_avalon_master_interface_0_avalon_master_0_read,          --                 .read
			avm_readdata      => sevensegment_avalon_master_interface_0_avalon_master_0_readdata,      --                 .readdata
			avm_write         => sevensegment_avalon_master_interface_0_avalon_master_0_write,         --                 .write
			avm_writedata     => sevensegment_avalon_master_interface_0_avalon_master_0_writedata,     --                 .writedata
			avm_waitrequest   => sevensegment_avalon_master_interface_0_avalon_master_0_waitrequest,   --                 .waitrequest
			avm_readdatavalid => sevensegment_avalon_master_interface_0_avalon_master_0_readdatavalid, --                 .readdatavalid
			rsi_reset_n       => rst_controller_reset_out_reset_ports_inv,                             --            reset.reset_n
			HEX7              => sevensegment_hex7,                                                    -- sevenseg_conduit.hex7
			HEX6              => sevensegment_hex6,                                                    --                 .hex6
			HEX5              => sevensegment_hex5,                                                    --                 .hex5
			HEX4              => sevensegment_hex4,                                                    --                 .hex4
			HEX3              => sevensegment_hex3,                                                    --                 .hex3
			HEX2              => sevensegment_hex2,                                                    --                 .hex2
			HEX1              => sevensegment_hex1,                                                    --                 .hex1
			HEX0              => sevensegment_hex0,                                                    --                 .hex0
			csi_clock         => sys_clk_clk                                                           --            clock.clk
		);

	mm_interconnect_1 : component EDAC_SDRAM_Controller_Demo_mm_interconnect_1
		port map (
			clk_0_clk_clk                                  => sys_clk_clk,                                                   --                                clk_0_clk.clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                -- nios2_gen2_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address               => nios2_gen2_0_data_master_address,                              --                 nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest           => nios2_gen2_0_data_master_waitrequest,                          --                                         .waitrequest
			nios2_gen2_0_data_master_byteenable            => nios2_gen2_0_data_master_byteenable,                           --                                         .byteenable
			nios2_gen2_0_data_master_read                  => nios2_gen2_0_data_master_read,                                 --                                         .read
			nios2_gen2_0_data_master_readdata              => nios2_gen2_0_data_master_readdata,                             --                                         .readdata
			nios2_gen2_0_data_master_write                 => nios2_gen2_0_data_master_write,                                --                                         .write
			nios2_gen2_0_data_master_writedata             => nios2_gen2_0_data_master_writedata,                            --                                         .writedata
			nios2_gen2_0_data_master_debugaccess           => nios2_gen2_0_data_master_debugaccess,                          --                                         .debugaccess
			nios2_gen2_0_instruction_master_address        => nios2_gen2_0_instruction_master_address,                       --          nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest    => nios2_gen2_0_instruction_master_waitrequest,                   --                                         .waitrequest
			nios2_gen2_0_instruction_master_read           => nios2_gen2_0_instruction_master_read,                          --                                         .read
			nios2_gen2_0_instruction_master_readdata       => nios2_gen2_0_instruction_master_readdata,                      --                                         .readdata
			edac_sdram_controller_0_porta_address          => mm_interconnect_1_edac_sdram_controller_0_porta_address,       --            edac_sdram_controller_0_porta.address
			edac_sdram_controller_0_porta_write            => mm_interconnect_1_edac_sdram_controller_0_porta_write,         --                                         .write
			edac_sdram_controller_0_porta_read             => mm_interconnect_1_edac_sdram_controller_0_porta_read,          --                                         .read
			edac_sdram_controller_0_porta_readdata         => mm_interconnect_1_edac_sdram_controller_0_porta_readdata,      --                                         .readdata
			edac_sdram_controller_0_porta_writedata        => mm_interconnect_1_edac_sdram_controller_0_porta_writedata,     --                                         .writedata
			edac_sdram_controller_0_porta_readdatavalid    => mm_interconnect_1_edac_sdram_controller_0_porta_readdatavalid, --                                         .readdatavalid
			edac_sdram_controller_0_porta_waitrequest      => mm_interconnect_1_edac_sdram_controller_0_porta_waitrequest,   --                                         .waitrequest
			nios2_gen2_0_debug_mem_slave_address           => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address,        --             nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write             => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write,          --                                         .write
			nios2_gen2_0_debug_mem_slave_read              => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read,           --                                         .read
			nios2_gen2_0_debug_mem_slave_readdata          => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata,       --                                         .readdata
			nios2_gen2_0_debug_mem_slave_writedata         => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata,      --                                         .writedata
			nios2_gen2_0_debug_mem_slave_byteenable        => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable,     --                                         .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest       => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest,    --                                         .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess       => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess,    --                                         .debugaccess
			onchip_memory2_0_s1_address                    => mm_interconnect_1_onchip_memory2_0_s1_address,                 --                      onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                      => mm_interconnect_1_onchip_memory2_0_s1_write,                   --                                         .write
			onchip_memory2_0_s1_readdata                   => mm_interconnect_1_onchip_memory2_0_s1_readdata,                --                                         .readdata
			onchip_memory2_0_s1_writedata                  => mm_interconnect_1_onchip_memory2_0_s1_writedata,               --                                         .writedata
			onchip_memory2_0_s1_byteenable                 => mm_interconnect_1_onchip_memory2_0_s1_byteenable,              --                                         .byteenable
			onchip_memory2_0_s1_chipselect                 => mm_interconnect_1_onchip_memory2_0_s1_chipselect,              --                                         .chipselect
			onchip_memory2_0_s1_clken                      => mm_interconnect_1_onchip_memory2_0_s1_clken,                   --                                         .clken
			onchip_memory2_0_s2_address                    => mm_interconnect_1_onchip_memory2_0_s2_address,                 --                      onchip_memory2_0_s2.address
			onchip_memory2_0_s2_write                      => mm_interconnect_1_onchip_memory2_0_s2_write,                   --                                         .write
			onchip_memory2_0_s2_readdata                   => mm_interconnect_1_onchip_memory2_0_s2_readdata,                --                                         .readdata
			onchip_memory2_0_s2_writedata                  => mm_interconnect_1_onchip_memory2_0_s2_writedata,               --                                         .writedata
			onchip_memory2_0_s2_byteenable                 => mm_interconnect_1_onchip_memory2_0_s2_byteenable,              --                                         .byteenable
			onchip_memory2_0_s2_chipselect                 => mm_interconnect_1_onchip_memory2_0_s2_chipselect,              --                                         .chipselect
			onchip_memory2_0_s2_clken                      => mm_interconnect_1_onchip_memory2_0_s2_clken                    --                                         .clken
		);

	irq_mapper : component EDAC_SDRAM_Controller_Demo_irq_mapper
		port map (
			clk        => sys_clk_clk,                    --       clk.clk
			reset      => rst_controller_reset_out_reset, -- clk_reset.reset
			sender_irq => nios2_gen2_0_irq_irq            --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => sys_rst_reset_n_ports_inv,          -- reset_in0.reset
			clk            => sys_clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	sys_rst_reset_n_ports_inv <= not sys_rst_reset_n;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of EDAC_SDRAM_Controller_Demo
